library verilog;
use verilog.vl_types.all;
entity MixColumn_vlg_vec_tst is
end MixColumn_vlg_vec_tst;
