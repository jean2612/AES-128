library verilog;
use verilog.vl_types.all;
entity MixColumn_vlg_check_tst is
    port(
        new_col_0       : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end MixColumn_vlg_check_tst;
